e866f14c59193e053e8ba5d38f4d55 ����   3 �  org/json/CDL  java/lang/Object <init> ()V Code
  	   LineNumberTable LocalVariableTable this Lorg/json/CDL; getValue *(Lorg/json/JSONTokener;)Ljava/lang/String; 
Exceptions  org/json/JSONException
    org/json/JSONTokener   next ()C  java/lang/StringBuffer
  	  java/lang/StringBuilder  Missing close quote '
  !  " (Ljava/lang/String;)V
  $ % & append (C)Ljava/lang/StringBuilder; ( '.
  * % + -(Ljava/lang/String;)Ljava/lang/StringBuilder;
  - . / toString ()Ljava/lang/String;
  1 2 3 syntaxError ,(Ljava/lang/String;)Lorg/json/JSONException;
  5 % 6 (C)Ljava/lang/StringBuffer;
  -
  9 :  back <  
  > ? @ nextTo (C)Ljava/lang/String; x Lorg/json/JSONTokener; c C q sb Ljava/lang/StringBuffer; StackMapTable rowToJSONArray ,(Lorg/json/JSONTokener;)Lorg/json/JSONArray; L org/json/JSONArray
 K 	
  O  
 K Q R S length ()I
 U Q V java/lang/String
 K X Y Z put ((Ljava/lang/Object;)Lorg/json/JSONArray; \ Bad character ' ^ ' (
  ` % a (I)Ljava/lang/StringBuilder; c ). ja Lorg/json/JSONArray; value Ljava/lang/String; rowToJSONObject A(Lorg/json/JSONArray;Lorg/json/JSONTokener;)Lorg/json/JSONObject;
  k I J
 K m n o toJSONObject +(Lorg/json/JSONArray;)Lorg/json/JSONObject; names r org/json/JSONObject rowToString ((Lorg/json/JSONArray;)Ljava/lang/String;
 K v w x opt (I)Ljava/lang/Object;
  -
 U { | } indexOf (I)I
 U  � � charAt (I)C
  � % � ,(Ljava/lang/String;)Ljava/lang/StringBuffer; i I object Ljava/lang/Object; string j toJSONArray ((Ljava/lang/String;)Lorg/json/JSONArray;
  !
  � � J
  � � � @(Lorg/json/JSONArray;Lorg/json/JSONTokener;)Lorg/json/JSONArray; <(Lorg/json/JSONArray;Ljava/lang/String;)Lorg/json/JSONArray;
  � h i jo Lorg/json/JSONObject;
 K � � � optJSONObject (I)Lorg/json/JSONObject;
 q � p � ()Lorg/json/JSONArray;
  � s t
 U � � � valueOf &(Ljava/lang/Object;)Ljava/lang/String;
  � . � <(Lorg/json/JSONArray;Lorg/json/JSONArray;)Ljava/lang/String;
 q � � � *(Lorg/json/JSONArray;)Lorg/json/JSONArray; 
SourceFile CDL.java !               /     *� �    
       .             
            H     �*� < ���	����    �          *   "   ,   '   ,   ,   {�=� Y� N*� <� � 6� 
� 	� *� Y�  � #'� )� ,� 0�-� 4W���-� 7�*� 8;�*� 8*,� =�    
   J    <  =  > < @ > C @ D H F M G R H U J e K  M � E � O � Q � R � T � U    *    � A B    � C D  @ M E D  H E F G  H    
 � ;� 	 �  	 I J          !     ~� KY� ML*� NM*� >,� +� P� ,� T� ,� �+,� WW,� ��� � 8
� � � +�*� Y[�  � #]� )� _b� )� ,� 0�*� >���    
   F    `  b  c  d  e * f , h 2 j 8 k ; m A n Q o S q f r r q v t { i    *    ~ A B    v d e   q f g   l C D  H    �  K� ! U" 	 h i           g     +� jM,� ,*� l� �    
   
    �  �          p e      A B    d e  H    �  K@ q 	 s t    �     ƻ Y� L=� �� 
+,� 4W*� uN-� �-� y:� T� {,� z� +
� z� !� z� � z� � ~"� I+"� 4W� T66� $� ~6 � "� 
+� 4W����+"� 4W� 
+� �W�*� P��V+
� 4W+� 7�    
   Z    �  �  �  �  �  � " � ( � : � N � b � i � p � v �  � � � � � � � � � � � � � � �    R    � d e    � F G  
 � � �   � � �  ( � � g  p 8 R �  s + � �    C D  H   ! 	�  
� I  U� � �  	 � �           6     � Y*� �� ��    
       �         � g   	 � J           3     	*� j*� ��    
       �        	 A B   	 � �           A     *� Y+� �� ��    
       �         p e      � g  	 � �           �     6*� 
*� P� �� KY� MM*+� �N-� � ,-� WW���,� P� �,�    
   .    �  �  �  �  �  � " � ( � + � 2 � 4 �    *    6 p e     6 A B   ! d e    � �  H    �  K�  q�  	 . t           �     /*� �L+� &+� �M,� � Y,� �� ��  ,*� �� )� ,��    
       �  � 
 �  �  � - �         / d e    ) � �    p e  H    � - q 	 . �           �     D*� 
*� P� �� Y� M>�  +� �:� ,*� �� �� �W�+� P���,� 7�    
   & 	       ! & 4 ?    4    D p e     D d e   / F G   ( � �  !  � �  H    �    �    �